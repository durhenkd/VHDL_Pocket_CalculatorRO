
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity ROM_COMENZI is
	 Port (CLK: in std_logic;
			 Adresa: in std_logic_vector(5 downto 0);
			 CS: in std_logic;
          D_ROM: out std_logic_vector(41 downto 0));
end ROM_COMENZI;

architecture Behavioral of ROM_COMENZI is

	signal adresa_temp: std_logic_vector(5 downto 0) := "000000";
	
begin
	
	process (CLK)
		begin
		if (rising_edge(CLK)) then
			if(CS = '0') then
				D_ROM <= "000000000000000000000000000000000000000000";
			else 
				case Adresa is 
	 when "000000" => D_ROM <= "000110011001010100000000000010100101000001";
	 when "000001" => D_ROM <= "000000000000000000000000000000000000000010";
	 when "000010" => D_ROM <= "100000000000000000000000000010000011000010";
	 when "000011" => D_ROM <= "000000000000000000001000000000000000000100";
	 when "000100" => D_ROM <= "000000100000000000000000000000000000000101";
	 when "000101" => D_ROM <= "000001000100000000000000000000000000000110";
	 when "000110" => D_ROM <= "001000000000000000000000000010000101000111";
	 when "000111" => D_ROM <= "000000000000101000000000000000000000001000";
	 when "001000" => D_ROM <= "100000000000000000000100000000001100001001";
	 when "001001" => D_ROM <= "100000000000000000000010000000010010001010";
	 when "001010" => D_ROM <= "100000000000000000000001000000010110001011";
	 when "001011" => D_ROM <= "100000000000000000000000100000100001000001";
	 when "001100" => D_ROM <= "000000000000000000000010101000000000001101";
	 when "001101" => D_ROM <= "000000000000000000000000000000000000001110";
	 when "001110" => D_ROM <= "000000000010000000000000000000000000001111";
	 when "001111" => D_ROM <= "000000000000000000000000000000010000010000";
	 when "010000" => D_ROM <= "100000000000000000000000010000010001111110";
	 when "010001" => D_ROM <= "000000000000000000000000000000000010111110";
	 when "010010" => D_ROM <= "000000000000000000000000000100000000010011";
	 when "010011" => D_ROM <= "000000000000000000000010100000000000010100";
	 when "010100" => D_ROM <= "000000000010000000000000000000000000010101";
	 when "010101" => D_ROM <= "000000000000000000000000000000010000111110";
	 when "010110" => D_ROM <= "000000000001000000000000000000000000010111";
	 when "010111" => D_ROM <= "000000000000000000000000000000001000011000";
	 when "011000" => D_ROM <= "000000000000000000010001010000000000011001";
	 when "011001" => D_ROM <= "000000000000000000000000001000000000011010";
	 when "011010" => D_ROM <= "000000000010000000000000000000000000011011";
	 when "011011" => D_ROM <= "000000000000000001000000000000000000011100";
	 when "011100" => D_ROM <= "000000000000000000000000000000001000011101";
	 when "011101" => D_ROM <= "100000000000000000000000000100011110011010";
	 when "011110" => D_ROM <= "000000000000000000000000000000010000011111";
	 when "011111" => D_ROM <= "100000000000000000000000010000100000111110";
	 when "100000" => D_ROM <= "000000000000000000000000000000000010111110";
	 when "100001" => D_ROM <= "100000000000000000000000001000100010100011";
	 when "100010" => D_ROM <= "000000000000000000000000000000000010111110";
	 when "100011" => D_ROM <= "000000000001000000010000000000001000100100";
	 when "100100" => D_ROM <= "000000000000000010000000000000000000100101";
	 when "100101" => D_ROM <= "000000000000000001000000000000000000100110";
	 when "100110" => D_ROM <= "000000000000000000000001100000000000100111";
	 when "100111" => D_ROM <= "000000000000000000000000000100000000101000";
	 when "101000" => D_ROM <= "000000000010000000000000000000000000101001";
	 when "101001" => D_ROM <= "000000000000000000000000000000001000101010";
	 when "101010" => D_ROM <= "100000000000000000000000000001101011101111";
	 when "101011" => D_ROM <= "000000000000000000010000000000000000101100";
	 when "101100" => D_ROM <= "000000000000000010000000000000000000101101";
	 when "101101" => D_ROM <= "000000000000000001000000000000000000101110";
	 when "101110" => D_ROM <= "000000000000000000000000001000000000110101";
	 when "101111" => D_ROM <= "010000000000000000100000000000000000110000";
	 when "110000" => D_ROM <= "000000000000100000000000000000000000110001";
	 when "110001" => D_ROM <= "000000000000000000010000000000000000110010";
	 when "110010" => D_ROM <= "000000000000000010000000000000000000110011";
	 when "110011" => D_ROM <= "000000000000000001000000000000000000110100";
	 when "110100" => D_ROM <= "000000000000000000000000000100000000110101";
	 when "110101" => D_ROM <= "000000000010000000000000000000000000110110";
	 when "110110" => D_ROM <= "000000000000000000000000000000001000110111";
	 when "110111" => D_ROM <= "100000000000000000000000000100111000101010";
	 when "111000" => D_ROM <= "100000000000000000000000000001111001111011";
	 when "111001" => D_ROM <= "000000000000000000000000001001000000111010";
	 when "111010" => D_ROM <= "000000000010000000000000000000000000111110";
	 when "111011" => D_ROM <= "010000000000000000100000000000000000111100";
	 when "111100" => D_ROM <= "000000000000100000000000000000000000111101";
	 when "111101" => D_ROM <= "000000000000000000000000000001000000111110";
	 when "111110" => D_ROM <= "000000000000000000000100000000010000111111";
	 when "111111" => D_ROM <= "000001100000000000000000000000000000000001";
	 when others => D_ROM <= "000000000000000000000000000000000000000000";
	 
	 end case;
	end if;
end if;

end process;
	
end Behavioral;

