
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity Screen_ROM is
	 Port (CLK: in std_logic;
			Adresa: in std_logic_vector(6 downto 0);
         CS: in std_logic;
          D_ROM: out std_logic_vector(20 downto 0) );
end Screen_ROM;

architecture Arh_Screen_ROM of Screen_ROM is

begin

process (CLK)
	begin
		if (rising_edge(CLK)) then
			if (CS = '0') then
				D_ROM <= "111111111111111111111";
			else
				case Adresa is
						when "0000000" => D_ROM <= "111111111111110000001";
						when "0000001" => D_ROM <= "111111111111111001111";
						when "0000010" => D_ROM <= "111111111111110010010";
						when "0000011" => D_ROM <= "111111111111110000110";
						when "0000100" => D_ROM <= "111111111111111001100";
						when "0000101" => D_ROM <= "111111111111110100100";
						when "0000110" => D_ROM <= "111111111111110100000";
						when "0000111" => D_ROM <= "111111111111110001111" ;
						when "0001000" => D_ROM <= "111111111111110000000";
						when "0001001" => D_ROM <= "111111111111110000100";
						when "0001010" => D_ROM <= "111111110011110000001";
	 when "0001011" => D_ROM <= "111111110011111001111";
	 when "0001100" => D_ROM <= "111111110011110010010";
	 when "0001101" => D_ROM <= "111111110011110000110";
	 when "0001110" => D_ROM <= "111111110011111001100";
	 when "0001111" => D_ROM <= "111111110011110100100";
	 when "0010000" => D_ROM <= "111111110011110100000";
	 when "0010001" => D_ROM <= "111111110011110001111";
	 when "0010010" => D_ROM <= "111111110011110000000";
	 when "0010011" => D_ROM <= "111111110011110000100";
	 when "0010100" => D_ROM <= "111111100100100000001";
	 when "0010101" => D_ROM <= "111111100100101001111";
	 when "0010110" => D_ROM <= "111111100100100010010";
	 when "0010111" => D_ROM <= "111111100100100000110";
	 when "0011000" => D_ROM <= "111111100100101001100";
	 when "0011001" => D_ROM <= "111111100100100100100";
	 when "0011010" => D_ROM <= "111111100100100100000";
	 when "0011011" => D_ROM <= "111111100100100001111";
	 when "0011100" => D_ROM <= "111111100100100000000";
	 when "0011101" => D_ROM <= "111111100100100000100";
	 when "0011110" => D_ROM <= "111111100001100000001";
	 when "0011111" => D_ROM <= "111111100001101001111";
	 when "0100000" => D_ROM <= "111111100001100010010";
	 when "0100001" => D_ROM <= "111111100001100000110";
	 when "0100010" => D_ROM <= "111111100001101001100";
	 when "0100011" => D_ROM <= "111111100001100100100";
	 when "0100100" => D_ROM <= "111111100001100100000";
	 when "0100101" => D_ROM <= "111111100001100001111";
	 when "0100110" => D_ROM <= "111111100001100000000";
	 when "0100111" => D_ROM <= "111111100001100000100";
	 when "0101000" => D_ROM <= "111111110011000000001";
	 when "0101001" => D_ROM <= "111111110011001001111";
	 when "0101010" => D_ROM <= "111111110011000010010";
	 when "0101011" => D_ROM <= "111111110011000000110";
	 when "0101100" => D_ROM <= "111111110011001001100";
	 when "0101101" => D_ROM <= "111111110011000100100";
	 when "0101110" => D_ROM <= "111111110011000100000";
	 when "0101111" => D_ROM <= "111111110011000001111";
	 when "0110000" => D_ROM <= "111111110011000000000";
	 when "0110001" => D_ROM <= "111111110011000000100";
	 when "0110010" => D_ROM <= "111111101001000000001";
	 when "0110011" => D_ROM <= "111111101001001001111";
	 when "0110100" => D_ROM <= "111111101001000010010";
	 when "0110101" => D_ROM <= "111111101001000000110";
	 when "0110110" => D_ROM <= "111111101001001001100";
	 when "0110111" => D_ROM <= "111111101001000100100";
	 when "0111000" => D_ROM <= "111111101001000100000";
	 when "0111001" => D_ROM <= "111111101001000001111";
	 when "0111010" => D_ROM <= "111111101001000000000";
	 when "0111011" => D_ROM <= "111111101001000000100";
	 when "0111100" => D_ROM <= "111111101000000000001";
	 when "0111101" => D_ROM <= "111111101000001001111";
	 when "0111110" => D_ROM <= "111111101000000010010";
	 when "0111111" => D_ROM <= "111111101000000000110";
	 when "1000000" => D_ROM <= "111111101000001001100";
	 when "1000001" => D_ROM <= "111111101000000100100";
	 when "1000010" => D_ROM <= "111111101000000100000";
	 when "1000011" => D_ROM <= "111111101000000001111";
	 when "1000100" => D_ROM <= "111111101000000000000";
	 when "1000101" => D_ROM <= "111111101000000000100";
	 when "1000110" => D_ROM <= "111111100011110000001";
	 when "1000111" => D_ROM <= "111111100011111001111";
	 when "1001000" => D_ROM <= "111111100011110010010";
	 when "1001001" => D_ROM <= "111111100011110000110";
	 when "1001010" => D_ROM <= "111111100011111001100";
	 when "1001011" => D_ROM <= "111111100011110100100";
	 when "1001100" => D_ROM <= "111111100011110100000";
	 when "1001101" => D_ROM <= "111111100011110001111";
	 when "1001110" => D_ROM <= "111111100011110000000";
	 when "1001111" => D_ROM <= "111111100011110000100";
	 when "1010000" => D_ROM <= "111111100000000000001";
	 when "1010001" => D_ROM <= "111111100000001001111";
	 when "1010010" => D_ROM <= "111111100000000010010";
	 when "1010011" => D_ROM <= "111111100000000000110";
	 when "1010100" => D_ROM <= "111111100000001001100";
	 when "1010101" => D_ROM <= "111111100000000100100";
	 when "1010110" => D_ROM <= "111111100000000100000";
	 when "1010111" => D_ROM <= "111111100000000001111";
	 when "1011000" => D_ROM <= "111111100000000000000";
	 when "1011001" => D_ROM <= "111111100000000000100";
	 when "1011010" => D_ROM <= "111111100001000000001";
	 when "1011011" => D_ROM <= "111111100001001001111";
	 when "1011100" => D_ROM <= "111111100001000010010";
	 when "1011101" => D_ROM <= "111111100001000000110";
	 when "1011110" => D_ROM <= "111111100001001001100";
	 when "1011111" => D_ROM <= "111111100001000100100";
	 when "1100000" => D_ROM <= "111111100001000100000";
	 when "1100001" => D_ROM <= "111111100001000001111";
	 when "1100010" => D_ROM <= "111111100001000000000";
	 when "1100011" => D_ROM <= "111111100001000000100";
	 when "1100100" => D_ROM <= "100111100000010000001";
	 when "1100101" => D_ROM <= "100111100000011001111";
	 when "1100110" => D_ROM <= "100111100000010010010";
	 when "1100111" => D_ROM <= "100111100000010000110";
	 when "1101000" => D_ROM <= "100111100000011001100";
	 when "1101001" => D_ROM <= "100111100000010100100";
	 when "1101010" => D_ROM <= "100111100000010100000";
	 when "1101011" => D_ROM <= "100111100000010001111";
	 when "1101100" => D_ROM <= "100111100000010000000";
	 when "1101101" => D_ROM <= "100111100000010000100";
	 when "1101110" => D_ROM <= "100111110011110000001";
	 when "1101111" => D_ROM <= "100111110011111001111";
	 when "1110000" => D_ROM <= "100111110011110010010";
	 when "1110001" => D_ROM <= "100111110011110000110";
	 when "1110010" => D_ROM <= "100111110011111001100";
	 when "1110011" => D_ROM <= "100111110011110100100";
	 when "1110100" => D_ROM <= "100111110011110100000";
	 when "1110101" => D_ROM <= "100111110011110001111";
	 when "1110110" => D_ROM <= "100111110011110000000";
	 when "1110111" => D_ROM <= "100111110011110000100";
	 when "1111000" => D_ROM <= "100111100100100000001";
	 when "1111001" => D_ROM <= "100111100100101001111";
	 when "1111010" => D_ROM <= "100111100100100010010";
	 when "1111011" => D_ROM <= "100111100100100000110";
	 when "1111100" => D_ROM <= "100111100100101001100";
	 when "1111101" => D_ROM <= "100111100100100100100";
	 when "1111110" => D_ROM <= "100111100100100100000";
	 when "1111111" => D_ROM <= "100111100100100001111";
	 when others => D_ROM <= "111111111111111111111";
	end case;
	end if;
	end if;
	end process;
end Arh_Screen_ROM;

